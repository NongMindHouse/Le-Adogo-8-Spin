`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:02:10 12/02/2023 
// Design Name: 
// Module Name:    header 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module header(horCnt,
				  verCnt,
				  clk,
				  rgbContent,
				  score,
				  endgamewin,
				  endgameLose
    );
	parameter headerStart = 31;
	parameter headerWidth = 4;
	parameter startSpr = 10;
	input [9:0] horCnt;
	input [9:0] verCnt;
	input clk;
	input [3:0] score;
	input endgamewin;
	input endgameLose;
	output reg [5:0] rgbContent = 0;
	reg [353:0] data_t = 354'b0;
	reg [9:0] magic = 0;
	
	always @(horCnt or verCnt) begin
		if(verCnt > headerStart && verCnt < headerStart+headerWidth) begin 
		//alphabet here
		
			rgbContent <= 6'b111111;
		end
		
		else if(verCnt < 32 && verCnt >= 0)
		      begin
		      if(horCnt >= (0+160) && horCnt < (354+160))
		      begin
		          if(endgamewin) begin 	
		          case(verCnt)
                  10'd00: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd01: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd02: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd03: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd04: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd05: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000011000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd06: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000011000000000000000001110000000000000110000000000000000000000000000000000000000000000000001100000000111100000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd07: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000011000000000000000011110000000000001110000000001100000000000000000000000000000000000000001100000011111100000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd08: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000011100000000000000111100000000000001110000000001100000000000000000000000000000000000000001110000011110000000000000000011000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd09: data_t = 354'b000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000001100000000000011110000000000000001100000000011100000000000000000000000110000000000000000110000000110000000111000000011000000000000000000000000000000000000011110001111110000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd10: data_t = 354'b000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000001100000000000011110000000000000001100000000011100000000000000000000000110000000000000000111000000110000000111000000011000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd11: data_t = 354'b000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000011100000000000000001111000000001111000000000000000001100000000011000000000000000000000000110000000000000000011000000110000000111110000011000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
                  10'd12: data_t = 354'b000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000011100000000000000001111100000111110000000000000000001100000000111000000000000000000000000110000000000000000011000000111000000111110000011100000000000000000000111000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000;
                  10'd13: data_t = 354'b000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000011110000000000000000011111111111000000000000000000001100000000111000000000000000000000000111000000000000000111000000011000000110111000001100000000000000000001111000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000;
                  10'd14: data_t = 354'b000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000011110001111000000000000111111100000000111111000000011100000001110000000000000000000000000011000000000000000110000000011000000111011100001100000000000000000011111000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd15: data_t = 354'b000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000011110011111000000000000000110000000011111111100000011100000001110000000000000000000000000011000000000000000110000000011000000111001110001100000000000000000011111000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd16: data_t = 354'b000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000011111111110000000000000001110000001111100001100000011000000001100000000000000000000000000111000000000000000110000000011000000011000110011100000000000000000111111000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd17: data_t = 354'b000000000000000000000000000000000000000000000000000000000111110000111100000000000000000000000011111111100000000000000001100000001111000001100000111000000001100000000000000000000000000110000001111000000110000000011000000011000111011000000000000000000111111000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd18: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000111111111100000000000000011100000001100000001100000111000000001100000000000000000000000000110000001111000000110000000011000000011000011111100000000011111111111111111000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd19: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000111111110000000000000000111000000001100000001100001110000000001100000000000000000000000000110000011111100000110000000011000000011000001111100000000011111111111111111110000000000111111011111000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd20: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000001111111110000000000000000110000000001100000001100001110000000011100000000000000000000000000111000011001110000110000000111000000011000001111110000000000111111111111111110000000000111000001111000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd21: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000001110000000001100000001100001100000000011100000000000000000000000000011000011000110000111000000110000000011000000011110000000000000111111111111100000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd22: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000011100000000001100000011100001100000000111000000000000000000000000000011000111000111000111000000110011100011100000001111000000000001111111111111000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd23: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011000000000001100000111100001100000000111000000000000000000000000000011000110000011100111000000110111100001100000000111000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd24: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000111000000000001111111110000001111111111110000000000000000000000000000011111110000001111110000000111110000001100000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd25: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000111000000000001111111110000001111111111110000000000000000000000000000011111110000000111100000000111100000001100000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd26: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000111100000000000110000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd27: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000011100000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd28: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd29: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd30: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd31: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  default: data_t = 354'b0;  
                  endcase;      
		          end
		          else if(endgameLose) begin 
		          case(verCnt)
                   10'd00: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd01: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd02: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd03: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd04: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000011000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd05: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111000000000000111100000000000000000000000000000000000000011111110000000000000000000000000111100000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd06: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001111000000000000111100000001110000000000000000000000000000111111111000000000000000000001111110000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd07: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000001111001111000000001111000000000000111110000011110000000000000000000000000001110000111100000000000000000001111100000000000000110011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd08: data_t = 354'b000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000111100000111000000001111100000000000110110000111110000000000000000000000000011110000011100000000000000000001100000001110000001110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd09: data_t = 354'b000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000111000000000000000001101110000000000110111001111110000001111111000000000000111000000001110000000000000000001100001111110000011100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd10: data_t = 354'b000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000001110000000000000000001100110000000000110011011100110000001111111000000000001110000000000110000000000000000001110111111000000011100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd11: data_t = 354'b000000000000000000000000000000000000000000000000000000000011111111111111100000000000001111110000000000001100000000000000000001100110000000000110011111000110000001100000000000000011100000000000110000000000000000000111111000000000111000000011000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd12: data_t = 354'b000000000000000000000000000000000000000000000000000000000011111111111111100000000000011111111000000000011100000000000000000011100111000000000110011110000110000001100000000000000011100000000000110000000000000000000111110000000001111110000111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd13: data_t = 354'b000000000000000000000000000000000000000000000000000000000001111111111111100000000000111111111000000000011100000000000000000011000011110000000110001110001110000011100000000000000011000000000000110000000000001100000111100000000001110111000111000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd14: data_t = 354'b000000000000000000000000000000000000000000000000000000000001111111111111100000000000111111111111100000111000000000011000000111011111110000000110001100001100000011000000000000000011000000000000110011000000011100000110000000000001100111111110000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd15: data_t = 354'b000000000000000000000000000000000000000000000000000000000000111111111111100000000000111111111111100000110000111111111000001111111111100000001110001100001100000011000000000000000011000000000000110011100000011000000110000111100011100011111100000000000111111100000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd16: data_t = 354'b000000000000000000000000000000000000000000000000000000000111000111111111100000000000111111111100000000110000111111111100001111110001100000001100000000011100000011110000000000000011000000000001110001100000111000000110001111100011000001110000000000001111111100000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd17: data_t = 354'b000000000000000000000000000000000000000000000000000000011111000011111111000000000000111111111000000000110000000000001100011111000001110000001100000000011000000111111111000000000011000000000001100001110000111000001110111100000111000000110000000000011111111110000000000011001111111100000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd18: data_t = 354'b000000000000000000000000000000000000000000000000000000011100001100011111000000000000111111111100000000110000000000001100111000000000110000011100000000111000001110111111000000000011000000000011100001111001110000001111111000000111000000110000000000011111111110000000000111001111111100000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd19: data_t = 354'b000000000000000000000000000000000000000000000000000000000000001100011000000000000000111110111100000000110000000000001101110000000000111000111000000000111000011100000000000000000011000000000011100000011101100000001111100000000110000000111000000000011111111110000000011111011111111100000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd20: data_t = 354'b000000000000000000000000000000000000000000000000000000000000111100011000000000000000000110001100000000111000000000011101100000000000111100110000000000110000011000000000000000000011100000001111000000011111100000001111000000000110000000111000000000011111111110000000011100111101111000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd21: data_t = 354'b000000000000000000000000000000000000000000000000000000000000111000111000000000000000001110000000000000011100000001111101100000000000011100110000000001110000011000000000000000000001110000111110000000001111100000001110000000000000000000011100000000011111111110000000000000111001100000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd22: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000111000000000000000001110000000000000001110000001110001100000000000001110110000000001110000011000000000000000000000111111111100000000000111100000000000000000000000000000011100000000000000000000000000000001111001100000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd23: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000001111111111100001100000000000001110000000000000000000111110000000000000000000111111110000000000000111000000000000000000000000000000000000000000000011001110000000000001110001100000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd24: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000011111111000001100000000000000110000000000000000000111111111110000000000000011111000000000000000011000000000000000000000000000000000000000000111011001111000000000001100011100000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd25: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011111110000000000000001110000000000000000000000000000000000000000000000000000000000001111011000111100000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd26: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110011000011100000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd27: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd28: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd29: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd30: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  10'd31: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                                  default: data_t = 354'b0;
                                  endcase;  		          
		          end
		          else begin 
		          case(verCnt)
                  10'd00: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd01: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
                  10'd02: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
                  10'd03: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000011110000010;
                  10'd04: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000011100000000000000000000000000000000000000000000000110000000000000001110000000000000000000000000000011110000000111111110000000000000000001110000000000111110000000000000000000000000000000000000000000000010000000011000000000000000000111010100110;
                  10'd05: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000111111100000000000000000000000000000000000000000000000110000000000000011110000011000000000000000000000111110000000111111110000000001100000011110000000001111111100000000000000001111111111110000000000000000111000000010000000000000000000001001111110;
                  10'd06: data_t = 354'b000000000000000000000011000000000000000000001111111111110000000000000000000011111000111100000000000000000011111111000000000000000000000000000000000000000000000000110000011000000111110000011100000000000011000001110110000000110000111100000001111111111100000000011100011100000000000000011111111111111100000000000000101000000010000000000000000000001001011010;
                  10'd07: data_t = 354'b000000000000000000000111000000000000000000011111111111111100000000000000000111100000000000000000000000000011100000000000111111111100000000000000000000000000000001110000011000000111111000001100000000000011000011110111000000110000011110000000111111111000000000011100011100000000000000111100000000011100000000000000101100111110011000111100000000011010000010;
                  10'd08: data_t = 354'b000000000000000000000111000000000000000000111100000000011100000000000000001111000000000000011111111110000011000000000000111111111100000000000000000000000000000001100000011000000110011000001100000000000011000111000011000000110000000110000000011000000000000000011000000000000000000001110000000000001100000000000001111100100110111000101101111000000000000000;
                  10'd09: data_t = 354'b000000000000000000001111000000000000000001110000000000001100000000000000001100000000000001111111111111100011100000000000110000001110000000000000000000000000000001100000011000001110011100001110000000001111000110000011100000111000000111000000011000000000000000011000000000000000000001110000000000001111000000000011000100101101101000101001001100000000000000;
                  10'd10: data_t = 354'b000000000000000000001111000000000000000001110000000000001111000000000000001100000000000001110000000111100001100000000000110000000111000000000000000000000000000001100000011000001100001100000110000000001110000110000001100000111000000011100000011000000000000000011000000000000000000011100000000000000111000000000010000100111101111000111001011111100000000000;
                  10'd11: data_t = 354'b000000000000000000001111100000000000000011100000000000000111000000000000001100000000000001100000000001100001100000000000110000000011000000000000000000000000000001100000011000011100001100000110000000111100011110000001100000011000000001100000011000000000000000011111000000000000000011000010000000100011000000000000000000000000000000001001110000000000000000;
                  10'd12: data_t = 354'b000000000000000000011111101111100000000011000011000001100011000000000000001110000000000001110000000001100001100000000000110000000011100000000000000000000000000001100000011100011000001110000110000000111000011100000001100000011000000001100000011000001110000000011111110000000000000011000011000001100011000000000000000000000000000000010000000000000000000000;
                  10'd13: data_t = 354'b000000000000000001111111111111100000000011000011000001100011000000000000000111100000000001110000000001100001100001110000110000000001100000000000000000000000000001100000001100111000000110000110000000110000111000000001110000011000000001100000011000011110000000000011110000000000000011000000000000000011000000000000000000001100000000100000000000000000000000;
                  10'd14: data_t = 354'b000000000000011111111111111111000000000011000000000000000011000000000000000011111100000000110000000001100001101111110000110000000001100000000000000000000000000001100000001110110000000110000110000000110000110000111111111000011000000001100000011100111100000000000000111110000000000011000000100010000011000000000000000000111110000000000000000000000000000000;
                  10'd15: data_t = 354'b000000000000011111111111111110000000000011000000111110000011000000000000000001111110000000110000000011100001111111100000110000001111100000000000000000000000000001100000000110110000000110000111000000110001111111111111111000011000000001100000001101110000000000000000011110000000000011000000110010000011000000000000000000111110000000000000000000000000000000;
                  10'd16: data_t = 354'b000000000000000111111111111100000000000011000000111110000011000000000000000000000111100000110000001111000011111100000000110111111111000000000000000000000000000001100000000111110000000110000011000001110001111111110000011000011000000001100000001111100000000000000000000110000000000011000000011110000011000000000000000111111110000000000000000000000000000000;
                  10'd17: data_t = 354'b000000000000000011111111111100000000000011000000011110000011000000000000000000000111110000110000111110000011000000000000110111111100000000000000000000000000000001100000000111100000000110000011100001100011100000000000011100011000000001100000001111000000000001100000000110000000000011100000000000000011000000001110000111111110000000000000000000000000000000;
                  10'd18: data_t = 354'b000000000000000001111111110000000000000011100000000000000011000000000000000000000000110000110000111000000011000000000000110011100000000000000000000000000000000001100000000111100000000110000011100001100011100000000000001100011000000001100000000110000000000001110000000110000000000001111111111111111111000000001111111111111110000000000000000000000000000000;
                  10'd19: data_t = 354'b000000000000000011111111100000000000000001111111111111111111000000000000000000000000110001111111110000000011000000000000110001110000000000000000000000000000000001100000000111100000000111000001100001100011000000000000001100011000000011100000000111000000000001111000000110000000000001111111111111111110000000000111111111111110000000000000000000000000000000;
                  10'd20: data_t = 354'b000000000000000011111111100000000000000001111111111111111110000000000000000000000000110001111111100000000111000000000000110000111000000000000000000000000000000001100000000111000000000011000001100011100011000000000000001100011100000011100000000011100000000000111000000110000000000000000000000000000000000000000011111111111111000000000000000000000000000000;
                  10'd21: data_t = 354'b000000000000000111111111110000000000000000000000000000000000000000110000000000000000110001110000000000000110000000000001110000011100000000000000000000000000000001100000001110000000000011000001100111000111000000000000001100001100000111000000000001100000000000011000000110000000000000000000000000000000000000000001111111111111100000000000000000000000000000;
                  10'd22: data_t = 354'b000000000000001111100011111000000000000000000000000000000000000000111000000000000000110001100000000000000110000000000001100000001111000000000000000000000000000001100000001110000000000011000001110110001110000000000000001110001110001111000000000001111000000000011100001110000000000001110000111000011110000000000011111111111111111000000000000000000000000000;
                  10'd23: data_t = 354'b000000000000011110000001111000000000000001110000111000011110000000111100000000000000110001100000000000000110000000000001100000000111000000000000000000000000000001100000001100000000000011000000111110001110000000000000000110001110011110000000000000111000000000001110011100000000000011110000111000011110000000000111111111111111111000000000000000000000000000;
                  10'd24: data_t = 354'b000000000000011000000000111100000000000011110000111000011110000000001110000000000001110001100000000000000110000001110001110000000011111000000000000000000000000001100000001100000000000011000000111100111100000000000000000000000111111100000000000000011111111100000111111000000000000011110001111000001111000000001111111111111110000000000000000000000000000000;
                  10'd25: data_t = 354'b000000000000011000000000111100000000000011110001111000001111000000000111000000000001110001100000000000000110000011110000110000000001111100000000000000000000000001100000001100000000000011000000111000111000000000000000000000000011110000000000000000011111111100000111111000000000000011100001111000001111000000011111111111111110000000000000000000000000000000;
                  10'd26: data_t = 354'b000000000000000000000000011100000000000011100001111000001111000000000011110000000111100001100000000000000110000111000000110000000000001110000000000000000000000001100000000000000000000000000000000000000000000000000000000000000011000000000000000000011100000000000011000000000000000011100001111000000111000000011100000000111110000000000000000000000000000000;
                  10'd27: data_t = 354'b000000000000000000000000000000000000000011100001111000000111000000000001111111111111000001100000000000000111111110000000110000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000;
                  10'd28: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000011111111110000001100000000000000111111100000000110000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000;
                  10'd29: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd30: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                  10'd31: data_t = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;		          
		           default: data_t = 354'b0;
		           endcase;
		          end
		         case(data_t[353-(horCnt-160)])
                      1: rgbContent <= 6'b111111;
                      0: rgbContent <= 6'b000000;
                      default: rgbContent <= 6'b000000;
                  endcase;
		      end
		      else 
                  rgbContent <= 6'b000000;               
	    end
	    else 
            rgbContent <= 6'b000000;
        end

endmodule