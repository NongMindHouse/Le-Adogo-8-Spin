`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:08:14 11/30/2023 
// Design Name: 
// Module Name:    drawPlayer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module drawPlayer(horCnt,
						verCnt,
						position,
						rgbContent
    );
	 input [9:0] horCnt;
	 input [9:0] verCnt;
	 input [9:0] position;
	 output reg [5:0] rgbContent = 6'bzzzzzz;
	 reg [32:0] data_t = 0;
	 
	always @(horCnt or verCnt or position) begin
			if(horCnt >= (position-15) && horCnt <= (position+15)) begin
				if(verCnt >= 416 && verCnt <= 447)begin
//fix here
                    case(verCnt - 416)
        10'd00: data_t = 33'b000000000000000000000000000000000;
        10'd01: data_t = 33'b000000000000000010000000000000000;
        10'd02: data_t = 33'b000000000000000010000000000000000;
        10'd03: data_t = 33'b000000000000000111000000000000000;
        10'd04: data_t = 33'b000000000000000101000000000000000;
        10'd05: data_t = 33'b000000000000000101000000000000000;
        10'd06: data_t = 33'b000000000000000101000000000000000;
        10'd07: data_t = 33'b000000100000000101000000001000000;
        10'd08: data_t = 33'b000000100000001111100000001000000;
        10'd09: data_t = 33'b000001110000011111110000011100000;
        10'd10: data_t = 33'b000001010000110000011000010100000;
        10'd11: data_t = 33'b000001010001100000011100010100000;
        10'd12: data_t = 33'b000001010011100011101110010100000;
        10'd13: data_t = 33'b000001010111100000011111010100000;
        10'd14: data_t = 33'b000001011111100000011111110100000;
        10'd15: data_t = 33'b000001011111110010011111110100000;
        10'd16: data_t = 33'b000001011111111111111111110100000;
        10'd17: data_t = 33'b000001111111111111111111111100000;
        10'd18: data_t = 33'b000011111111111111111111111110000;
        10'd19: data_t = 33'b000111111111111111111111111111000;
        10'd20: data_t = 33'b000111111111111111111111111111000;
        10'd21: data_t = 33'b001111111111111111111111111111100;
        10'd22: data_t = 33'b001111111111111111111111111111100;
        10'd23: data_t = 33'b011111111100011111110001111111110;
        10'd24: data_t = 33'b011111111000001111100000111111110;
        10'd25: data_t = 33'b011111110000111111111000011111110;
        10'd26: data_t = 33'b011111100001111111111100001111110;
        10'd27: data_t = 33'b011111000000000000000000000111110;
        10'd28: data_t = 33'b001110000000000000000000000011100;
        10'd29: data_t = 33'b000000000000000000000000000000000;
        10'd30: data_t = 33'b000000000000000000000000000000000;
        10'd31: data_t = 33'b000000000000000000000000000000000;
        10'd32: data_t = 33'b000000000000000000000000000000000;
        default: data_t = 33'b000000000000000000000000000000000;        
                endcase
                
                case(data_t[horCnt-(position-16)])
                    1: rgbContent <= 6'b111111;
                    0: rgbContent <= 6'b000000;
                    default: rgbContent <= 6'b000000;
                endcase
            end
			else 
                rgbContent = 6'b000000;            
            end
 //fix here
			else 
				rgbContent = 6'b000000;
	        end

endmodule
